module rxv

import time

pub interface Duration {
	duration() time.Duration
}
