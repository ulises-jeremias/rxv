module rxv
