module rxv

struct ChannelIterable {
}
