module rxv

import context
import sync

type OperatorFactoryFn = fn () Operator
